module UART_transmitter
      #(parameter D_BIT = 8, 
		            SB_TICK = 16
		)
		(
		input clk, rst,
		input tx_start, s_tick,
		input [D_BIT-1:0] d_in,
		output wire tx,
		output reg tx_done_tick
		);
		
localparam [1:0] 
         idle = 2'b00, 
			start = 2'b01, 
			data = 2'b10, 
			stop = 2'b11;	
			
reg [1:0] state_reg, state_next;	
reg [3:0] s_reg, s_next;         
reg [2:0] n_reg, n_next;
reg [D_BIT-1:0] b_reg, b_next;
reg tx_reg, tx_next;

always@(posedge clk, posedge rst)
begin
     if(rst)
	  begin
	     state_reg <= idle;
		  s_reg <= 0;
		  n_reg <= 0;
		  b_reg <= 0;
		  tx_reg <= 1'b1;
	  end
	  else
	  begin 
	     state_reg <= state_next;
		  s_reg <= s_next;
		  n_reg <= n_next;
		  b_reg <= b_next;
		  tx_reg <= tx_next;
	  end  
end
always @*
begin
     state_next <= state_reg;
	  s_next <= s_reg;
	  n_next <= n_reg;
	  b_next <= b_reg;
	  tx_next <= tx_reg;
	  tx_done_tick <= 1'b0;
     case(state_reg)
	       idle:  begin
			         tx_next = 1'b1;
			        if(tx_start == 0)
					  begin
					     state_next = start;
						  s_next = 0;
						  b_next = d_in;
					  end
					  end
		    start: begin
			        tx_next = 1'b0;
			 		  if(s_tick == 1'b1)
			           if(s_reg == 4'd15)
						     begin
						     s_next = 0;
							  n_next = 0;
							  state_next = data;
							  end
						  else 
					        s_next = s_reg + 1;
					  end
			 data: begin
			       tx_next = b_reg[0];
			       if(s_tick == 1'b1)
					     if(s_reg == 4'd15)
						  begin
						     s_next = 0;
							  b_next = b_reg >> 1;
							  if(n_reg == (D_BIT - 1))
							    state_next = stop;
							  else 
							    n_next = n_reg + 1;
						  end
						  else 
						      s_next = s_reg + 1;
				 	end
	       stop: begin
			       tx_next = 1'b0;
			       if(s_tick == 1'b1)
					    if(s_reg == (SB_TICK - 1))
						     begin
							  tx_done_tick = 1'b1;
							  state_next = idle;
							  end
						 else 
							  s_next = s_reg + 1;		 					 
                end    
	  endcase
end
assign tx = tx_reg;

endmodule 
				
	   
